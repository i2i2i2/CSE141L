/*****************************************************************************
  File Name:    ALU.sv
  Author:       Chenxu Jiang
                DingCheng Hu
  Date:         Apr 29, 2017
  Description:  ALU
                Input   
*****************************************************************************/
