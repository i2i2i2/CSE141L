/*****************************************************************************
  File Name:    InstrDecoder.sv
  Author:       Chenxu Jiang
                DingCheng Hu
  Date:         Apr 29, 2017
  Description:  decode instruction, control state of all units
                TBD
*****************************************************************************/
