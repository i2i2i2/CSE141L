/*****************************************************************************
  File Name:    SingleCycleCPU.sv
  Author:       Chenxu Jiang
                DingCheng Hu
  Date:         Apr 29, 2017
  Description:  put every module together
*****************************************************************************/
`timescale 1s / 1s
`include "ALU.sv"
`include "dataMem.sv"
`include "InstrFetch.sv"
`include "InstrDecoder.sv"
`include "RegsFile.sv"

module SingleCycleCPU;

  wire[8:0]     instr, control;
  wire[7:0]     regData, addr, dataIn, dataOut, result, srcA, srcB, srcC;
  wire[2:0]     read1, read2, writeReg, regSrc;
  wire[1:0]     branchCtrl;
  wire          memOp, writeBranch, isReg1, isReg2, isReg3, isWrite, writeFlip,
                isRegW, writeFlag, flag0, flag1, flip0, flip2, branchResult, halt;

  reg           init, CLK;

  InstrFetch IF(init, halt, writeBranch, branchResult, branchCtrl, CLK, instr);
  InstrDecode ID(instr, writeBranch, branchCtrl, halt, control, read1, isReg1,
      read2, isReg2, isReg3, isWrite, writeReg, isRegW, regData, writeFlip,
      writeFlag, memOp, regSrc);
  RegsFile RF(read1, isReg1, read2, isReg2, isReg3, isWrite, writeReg,
      result, regData, dataOut, srcA, regSrc, isRegW, flip0, writeFlip,
      flag0, writeFlip, CLK, srcA, srcB, srcC, flip1, flag1);
  ALU ALU0(srcA, srcB, srcC, flag1, flip1, control, result, flag0, flip0, branchResult);
  dataMem M(srcA, srcB, memOp, CLK, dataOut);

  always begin
    #1 CLK = 1;
    #1 CLK = 0;
  end

  initial begin
    $dumpfile("CPU.vcd");
    $dumpvars(0, SingleCycleCPU);

    $monitor ("%b:  %b", CLK, instr);
    init = 1'b1;
    #2 init = 1'b0;
  end

  initial begin
    #500 $finish;
  end

endmodule
